

// 
// Module: tb
// 
// Notes:
// - Top level simulation testbench.
//

//`timescale 1ns/1ns
//`define WAVES_FILE "./work/waves-rx.vcd"

module tb();
    
reg        clk          ; // Top level system clock input.
reg rst;
reg neg_clk; 
reg neg_rst ; 
reg        resetn       ;
reg        uart_rxd     ; // UART Recieve pin.

reg        uart_rx_en   ; // Recieve enable
//wire [8:0] res;
wire       uart_rx_break; // Did we get a BREAK message?
wire       uart_rx_valid; // Valid data recieved and available.
wire [7:0] uart_rx_data ; // The recieved data.
wire [31:0] inst ; 
wire [31:0] inst_mem ; 

reg rst_pin ; 
wire write_done ; 


// Bit rate of the UART line we are testing.
localparam BIT_RATE = 9600;
localparam BIT_P    = (1000000000/BIT_RATE);


// Period and frequency of the system clock.
localparam CLK_HZ   = 50000000;
localparam CLK_P    = 1000000000/ CLK_HZ;

reg slow_clk = 0;


// Make the clock tick.
always begin #(CLK_P/2) clk  = ~clk; end   
always begin #(CLK_P/2) neg_clk  = ~neg_clk; end     
always begin #(CLK_P*2) slow_clk <= !slow_clk;end



task write_instruction;
    input [31:0] instruction;
    begin
            @(posedge clk);
            send_byte(instruction[7:0]);
            check_byte(instruction[7:0]);
            @(posedge clk);
            send_byte(instruction[15:8]);
            check_byte(instruction[15:8]);
            
            @(posedge clk);
            send_byte(instruction[23:16]);
            check_byte(instruction[23:16]);
            
            @(posedge clk);
            send_byte(instruction[31:24]);
            check_byte(instruction[31:24]);
    end
    endtask

task send_byte;
    input [7:0] to_send;
    integer i;
    begin


        #BIT_P;  uart_rxd = 1'b0;
        for(i=0; i < 8; i = i+1) begin
            #BIT_P;  uart_rxd = to_send[i];
        end
        #BIT_P;  uart_rxd = 1'b1;
        #1000;
    end
endtask


// Checks that the output of the UART is the value we expect.
integer passes = 0;
integer fails  = 0;
task check_byte;
    input [7:0] expected_value;
    begin
        if(uart_rx_data == expected_value) begin
            passes = passes + 1;
            $display("%d/%d/%d [PASS] Expected %b and got %b", 
                     passes,fails,passes+fails,
                     expected_value, uart_rx_data);
        end else begin
            fails  = fails  + 1;
            $display("%d/%d/%d [FAIL] Expected %b and got %b", 
                     passes,fails,passes+fails,
                     expected_value, uart_rx_data);
        end
    end
endtask


initial 
begin 
    $dumpfile("waveform.vcd");
    $dumpvars(0,tb);
end 

reg [7:0] input_wires; 
wire [31:8] output_wires ; 
wire [2:0] pc ; 


reg [7:0] to_send;
initial begin
    rst=1;
    rst_pin=1; 
    neg_rst = 1; 
    resetn  = 1'b0;
    clk     = 1'b0;
    neg_clk = 1; 
    neg_rst = ~clk ;
    uart_rxd = 1'b1;
    neg_clk = 1'b1; 
    input_wires = 8'b00010001;
    #4000
    resetn = 1'b1;
    rst=0;
    neg_rst = 0; 
    rst_pin = 0 ; 
  

    uart_rx_en = 1'b1;
    @(posedge slow_clk);write_instruction(32'h00000000); 
    @(posedge slow_clk);write_instruction(32'h00000000); 
    @(posedge slow_clk);write_instruction(32'hfd010113); 
    @(posedge slow_clk);write_instruction(32'h02812623); 
    @(posedge slow_clk);write_instruction(32'h03010413); 
    @(posedge slow_clk);write_instruction(32'hfca42e23); 
    @(posedge slow_clk);write_instruction(32'hfdc42783); 
    @(posedge slow_clk);write_instruction(32'h00100713); 
    @(posedge slow_clk);write_instruction(32'h00f717b3); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00ff6f33); 
    @(posedge slow_clk);write_instruction(32'h00000013); 
    @(posedge slow_clk);write_instruction(32'h02c12403); 
    @(posedge slow_clk);write_instruction(32'h03010113); 
    @(posedge slow_clk);write_instruction(32'h00008067); 
    @(posedge slow_clk);write_instruction(32'hfd010113); 
    @(posedge slow_clk);write_instruction(32'h02812623); 
    @(posedge slow_clk);write_instruction(32'h03010413); 
    @(posedge slow_clk);write_instruction(32'hfca42e23); 
    @(posedge slow_clk);write_instruction(32'hfdc42783); 
    @(posedge slow_clk);write_instruction(32'h00100713); 
    @(posedge slow_clk);write_instruction(32'h00f717b3); 
    @(posedge slow_clk);write_instruction(32'hfff7c793); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00ff7f33); 
    @(posedge slow_clk);write_instruction(32'h00000013); 
    @(posedge slow_clk);write_instruction(32'h02c12403); 
    @(posedge slow_clk);write_instruction(32'h03010113); 
    @(posedge slow_clk);write_instruction(32'h00008067); 
    @(posedge slow_clk);write_instruction(32'hfd010113); 
    @(posedge slow_clk);write_instruction(32'h02812623); 
    @(posedge slow_clk);write_instruction(32'h03010413); 
    @(posedge slow_clk);write_instruction(32'hfca42e23); 
    @(posedge slow_clk);write_instruction(32'hfe042623); 
    @(posedge slow_clk);write_instruction(32'h000f0793); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'hfdc42783); 
    @(posedge slow_clk);write_instruction(32'hfec42703); 
    @(posedge slow_clk);write_instruction(32'h40f757b3); 
    @(posedge slow_clk);write_instruction(32'h0017f793); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'h02c12403); 
    @(posedge slow_clk);write_instruction(32'h03010113); 
    @(posedge slow_clk);write_instruction(32'h00008067); 
    @(posedge slow_clk);write_instruction(32'hfe010113); 
    @(posedge slow_clk);write_instruction(32'h00112e23); 
    @(posedge slow_clk);write_instruction(32'h00812c23); 
    @(posedge slow_clk);write_instruction(32'h02010413); 
    @(posedge slow_clk);write_instruction(32'hfea42623); 
    @(posedge slow_clk);write_instruction(32'hfeb42423); 
    @(posedge slow_clk);write_instruction(32'hfec42223); 
    @(posedge slow_clk);write_instruction(32'hfed42023); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h0007a023); 
    @(posedge slow_clk);write_instruction(32'hfe842503); 
    @(posedge slow_clk);write_instruction(32'hf5dff0ef); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'hf1dff0ef); 
    @(posedge slow_clk);write_instruction(32'hfe042783); 
    @(posedge slow_clk);write_instruction(32'h00100713); 
    @(posedge slow_clk);write_instruction(32'h00e7a023); 
    @(posedge slow_clk);write_instruction(32'h00000013); 
    @(posedge slow_clk);write_instruction(32'h01c12083); 
    @(posedge slow_clk);write_instruction(32'h01812403); 
    @(posedge slow_clk);write_instruction(32'h02010113); 
    @(posedge slow_clk);write_instruction(32'h00008067); 
    @(posedge slow_clk);write_instruction(32'hfe010113); 
    @(posedge slow_clk);write_instruction(32'h00112e23); 
    @(posedge slow_clk);write_instruction(32'h00812c23); 
    @(posedge slow_clk);write_instruction(32'h02010413); 
    @(posedge slow_clk);write_instruction(32'hfea42623); 
    @(posedge slow_clk);write_instruction(32'hfeb42423); 
    @(posedge slow_clk);write_instruction(32'hfec42223); 
    @(posedge slow_clk);write_instruction(32'hfed42023); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h0007a023); 
    @(posedge slow_clk);write_instruction(32'hfe842503); 
    @(posedge slow_clk);write_instruction(32'hf05ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'hec5ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfe042783); 
    @(posedge slow_clk);write_instruction(32'h00100713); 
    @(posedge slow_clk);write_instruction(32'h00e7a023); 
    @(posedge slow_clk);write_instruction(32'h00000013); 
    @(posedge slow_clk);write_instruction(32'h01c12083); 
    @(posedge slow_clk);write_instruction(32'h01812403); 
    @(posedge slow_clk);write_instruction(32'h02010113); 
    @(posedge slow_clk);write_instruction(32'h00008067); 
    @(posedge slow_clk);write_instruction(32'hfd010113); 
    @(posedge slow_clk);write_instruction(32'h02112623); 
    @(posedge slow_clk);write_instruction(32'h02812423); 
    @(posedge slow_clk);write_instruction(32'h03010413); 
    @(posedge slow_clk);write_instruction(32'hfca42e23); 
    @(posedge slow_clk);write_instruction(32'hfcb42c23); 
    @(posedge slow_clk);write_instruction(32'hfcc42a23); 
    @(posedge slow_clk);write_instruction(32'hfe042623); 
    @(posedge slow_clk);write_instruction(32'hfd442503); 
    @(posedge slow_clk);write_instruction(32'heb5ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfd842503); 
    @(posedge slow_clk);write_instruction(32'he75ff0ef); 
    @(posedge slow_clk);write_instruction(32'h0100006f); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00178793); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'hfec42703); 
    @(posedge slow_clk);write_instruction(32'h3e800793); 
    @(posedge slow_clk);write_instruction(32'hfef716e3); 
    @(posedge slow_clk);write_instruction(32'hfd842503); 
    @(posedge slow_clk);write_instruction(32'he89ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'he49ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00000013); 
    @(posedge slow_clk);write_instruction(32'h02c12083); 
    @(posedge slow_clk);write_instruction(32'h02812403); 
    @(posedge slow_clk);write_instruction(32'h03010113); 
    @(posedge slow_clk);write_instruction(32'h00008067); 
    @(posedge slow_clk);write_instruction(32'hf9010113); 
    @(posedge slow_clk);write_instruction(32'h06112623); 
    @(posedge slow_clk);write_instruction(32'h06812423); 
    @(posedge slow_clk);write_instruction(32'h07010413); 
    @(posedge slow_clk);write_instruction(32'hfca42e23); 
    @(posedge slow_clk);write_instruction(32'hfcb42c23); 
    @(posedge slow_clk);write_instruction(32'hfcc42a23); 
    @(posedge slow_clk);write_instruction(32'hfcd42823); 
    @(posedge slow_clk);write_instruction(32'hfce42623); 
    @(posedge slow_clk);write_instruction(32'hfcf42423); 
    @(posedge slow_clk);write_instruction(32'hfd042223); 
    @(posedge slow_clk);write_instruction(32'hfd142023); 
    @(posedge slow_clk);write_instruction(32'h00f00793); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'h02d00793); 
    @(posedge slow_clk);write_instruction(32'hfef42423); 
    @(posedge slow_clk);write_instruction(32'hfe042223); 
    @(posedge slow_clk);write_instruction(32'hfe042023); 
    @(posedge slow_clk);write_instruction(32'hfe040793); 
    @(posedge slow_clk);write_instruction(32'h02f12623); 
    @(posedge slow_clk);write_instruction(32'hfe440793); 
    @(posedge slow_clk);write_instruction(32'h02f12423); 
    @(posedge slow_clk);write_instruction(32'h02012223); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h02f12023); 
    @(posedge slow_clk);write_instruction(32'h01c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'h01842783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'h01442783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'h01042783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'h00c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'h00842783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'h00442783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'h00042783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfc042883); 
    @(posedge slow_clk);write_instruction(32'hfc442803); 
    @(posedge slow_clk);write_instruction(32'hfc842783); 
    @(posedge slow_clk);write_instruction(32'hfcc42703); 
    @(posedge slow_clk);write_instruction(32'hfd042683); 
    @(posedge slow_clk);write_instruction(32'hfd442603); 
    @(posedge slow_clk);write_instruction(32'hfd842583); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'h09c000ef); 
    @(posedge slow_clk);write_instruction(32'hfe040793); 
    @(posedge slow_clk);write_instruction(32'h02f12623); 
    @(posedge slow_clk);write_instruction(32'hfe440793); 
    @(posedge slow_clk);write_instruction(32'h02f12423); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f12223); 
    @(posedge slow_clk);write_instruction(32'hfe842783); 
    @(posedge slow_clk);write_instruction(32'h02f12023); 
    @(posedge slow_clk);write_instruction(32'h01c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'h01842783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'h01442783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'h01042783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'h00c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'h00842783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'h00442783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'h00042783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfc042883); 
    @(posedge slow_clk);write_instruction(32'hfc442803); 
    @(posedge slow_clk);write_instruction(32'hfc842783); 
    @(posedge slow_clk);write_instruction(32'hfcc42703); 
    @(posedge slow_clk);write_instruction(32'hfd042683); 
    @(posedge slow_clk);write_instruction(32'hfd442603); 
    @(posedge slow_clk);write_instruction(32'hfd842583); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'h018000ef); 
    @(posedge slow_clk);write_instruction(32'h00000013); 
    @(posedge slow_clk);write_instruction(32'h06c12083); 
    @(posedge slow_clk);write_instruction(32'h06812403); 
    @(posedge slow_clk);write_instruction(32'h07010113); 
    @(posedge slow_clk);write_instruction(32'h00008067); 
    @(posedge slow_clk);write_instruction(32'hfa010113); 
    @(posedge slow_clk);write_instruction(32'h04112e23); 
    @(posedge slow_clk);write_instruction(32'h04812c23); 
    @(posedge slow_clk);write_instruction(32'h06010413); 
    @(posedge slow_clk);write_instruction(32'hfaa42e23); 
    @(posedge slow_clk);write_instruction(32'hfab42c23); 
    @(posedge slow_clk);write_instruction(32'hfac42a23); 
    @(posedge slow_clk);write_instruction(32'hfad42823); 
    @(posedge slow_clk);write_instruction(32'hfae42623); 
    @(posedge slow_clk);write_instruction(32'hfaf42423); 
    @(posedge slow_clk);write_instruction(32'hfb042223); 
    @(posedge slow_clk);write_instruction(32'hfb142023); 
    @(posedge slow_clk);write_instruction(32'hfe042623); 
    @(posedge slow_clk);write_instruction(32'hfe042423); 
    @(posedge slow_clk);write_instruction(32'hfe042223); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hfcf42c23); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hfcf42a23); 
    @(posedge slow_clk);write_instruction(32'hfc042823); 
    @(posedge slow_clk);write_instruction(32'hfc042623); 
    @(posedge slow_clk);write_instruction(32'hfc042423); 
    @(posedge slow_clk);write_instruction(32'hfc042223); 
    @(posedge slow_clk);write_instruction(32'hfe042023); 
    @(posedge slow_clk);write_instruction(32'hfc042e23); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h00078c63); 
    @(posedge slow_clk);write_instruction(32'h02842783); 
    @(posedge slow_clk);write_instruction(32'h00078863); 
    @(posedge slow_clk);write_instruction(32'hfc042c23); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hfcf42823); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h00078c63); 
    @(posedge slow_clk);write_instruction(32'h02c42783); 
    @(posedge slow_clk);write_instruction(32'h00078863); 
    @(posedge slow_clk);write_instruction(32'hfc042a23); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hfcf42623); 
    @(posedge slow_clk);write_instruction(32'h02442703); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f71a63); 
    @(posedge slow_clk);write_instruction(32'hfbc42503); 
    @(posedge slow_clk);write_instruction(32'hc99ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02078263); 
    @(posedge slow_clk);write_instruction(32'hfd040713); 
    @(posedge slow_clk);write_instruction(32'hfd840793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'h01042603); 
    @(posedge slow_clk);write_instruction(32'hfac42583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'hd09ff0ef); 
    @(posedge slow_clk);write_instruction(32'h0380006f); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h02079863); 
    @(posedge slow_clk);write_instruction(32'hfb842503); 
    @(posedge slow_clk);write_instruction(32'hc61ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02078063); 
    @(posedge slow_clk);write_instruction(32'hfd040713); 
    @(posedge slow_clk);write_instruction(32'hfd840793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'h01842603); 
    @(posedge slow_clk);write_instruction(32'hfa442583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'hcd1ff0ef); 
    @(posedge slow_clk);write_instruction(32'h02442703); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f71a63); 
    @(posedge slow_clk);write_instruction(32'hfb442503); 
    @(posedge slow_clk);write_instruction(32'hc29ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02078263); 
    @(posedge slow_clk);write_instruction(32'hfcc40713); 
    @(posedge slow_clk);write_instruction(32'hfd440793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'h01442603); 
    @(posedge slow_clk);write_instruction(32'hfa842583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'hc99ff0ef); 
    @(posedge slow_clk);write_instruction(32'h0380006f); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h38079463); 
    @(posedge slow_clk);write_instruction(32'hfb042503); 
    @(posedge slow_clk);write_instruction(32'hbf1ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h36078c63); 
    @(posedge slow_clk);write_instruction(32'hfcc40713); 
    @(posedge slow_clk);write_instruction(32'hfd440793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'h01c42603); 
    @(posedge slow_clk);write_instruction(32'hfa042583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'hc61ff0ef); 
    @(posedge slow_clk);write_instruction(32'h3580006f); 
    @(posedge slow_clk);write_instruction(32'hfd042783); 
    @(posedge slow_clk);write_instruction(32'h06078663); 
    @(posedge slow_clk);write_instruction(32'h02442703); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h06f71063); 
    @(posedge slow_clk);write_instruction(32'hfbc42503); 
    @(posedge slow_clk);write_instruction(32'hbadff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050713); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f70663); 
    @(posedge slow_clk);write_instruction(32'h02042703); 
    @(posedge slow_clk);write_instruction(32'h00070793); 
    @(posedge slow_clk);write_instruction(32'h00579793); 
    @(posedge slow_clk);write_instruction(32'h40e787b3); 
    @(posedge slow_clk);write_instruction(32'h00279793); 
    @(posedge slow_clk);write_instruction(32'h00e787b3); 
    @(posedge slow_clk);write_instruction(32'h00379793); 
    @(posedge slow_clk);write_instruction(32'h00078713); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h02e7c263); 
    @(posedge slow_clk);write_instruction(32'hfc840713); 
    @(posedge slow_clk);write_instruction(32'hfd040793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'h00042603); 
    @(posedge slow_clk);write_instruction(32'h01042583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'hb99ff0ef); 
    @(posedge slow_clk);write_instruction(32'h06c0006f); 
    @(posedge slow_clk);write_instruction(32'hfd042783); 
    @(posedge slow_clk);write_instruction(32'h06078263); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h04079e63); 
    @(posedge slow_clk);write_instruction(32'hfb842503); 
    @(posedge slow_clk);write_instruction(32'hb41ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050713); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f70663); 
    @(posedge slow_clk);write_instruction(32'h02042703); 
    @(posedge slow_clk);write_instruction(32'h00070793); 
    @(posedge slow_clk);write_instruction(32'h00579793); 
    @(posedge slow_clk);write_instruction(32'h40e787b3); 
    @(posedge slow_clk);write_instruction(32'h00279793); 
    @(posedge slow_clk);write_instruction(32'h00e787b3); 
    @(posedge slow_clk);write_instruction(32'h00379793); 
    @(posedge slow_clk);write_instruction(32'h00078713); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h02e7c063); 
    @(posedge slow_clk);write_instruction(32'hfc840713); 
    @(posedge slow_clk);write_instruction(32'hfd040793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'h00842603); 
    @(posedge slow_clk);write_instruction(32'h01842583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'hb2dff0ef); 
    @(posedge slow_clk);write_instruction(32'hfcc42783); 
    @(posedge slow_clk);write_instruction(32'h06078663); 
    @(posedge slow_clk);write_instruction(32'h02442703); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h06f71063); 
    @(posedge slow_clk);write_instruction(32'hfb442503); 
    @(posedge slow_clk);write_instruction(32'had5ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050713); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f70663); 
    @(posedge slow_clk);write_instruction(32'h02042703); 
    @(posedge slow_clk);write_instruction(32'h00070793); 
    @(posedge slow_clk);write_instruction(32'h00579793); 
    @(posedge slow_clk);write_instruction(32'h40e787b3); 
    @(posedge slow_clk);write_instruction(32'h00279793); 
    @(posedge slow_clk);write_instruction(32'h00e787b3); 
    @(posedge slow_clk);write_instruction(32'h00379793); 
    @(posedge slow_clk);write_instruction(32'h00078713); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h02e7c263); 
    @(posedge slow_clk);write_instruction(32'hfc440713); 
    @(posedge slow_clk);write_instruction(32'hfcc40793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'h00442603); 
    @(posedge slow_clk);write_instruction(32'h01442583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'hac1ff0ef); 
    @(posedge slow_clk);write_instruction(32'h06c0006f); 
    @(posedge slow_clk);write_instruction(32'hfcc42783); 
    @(posedge slow_clk);write_instruction(32'h06078263); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h04079e63); 
    @(posedge slow_clk);write_instruction(32'hfb042503); 
    @(posedge slow_clk);write_instruction(32'ha69ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050713); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f70663); 
    @(posedge slow_clk);write_instruction(32'h02042703); 
    @(posedge slow_clk);write_instruction(32'h00070793); 
    @(posedge slow_clk);write_instruction(32'h00579793); 
    @(posedge slow_clk);write_instruction(32'h40e787b3); 
    @(posedge slow_clk);write_instruction(32'h00279793); 
    @(posedge slow_clk);write_instruction(32'h00e787b3); 
    @(posedge slow_clk);write_instruction(32'h00379793); 
    @(posedge slow_clk);write_instruction(32'h00078713); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h02e7c063); 
    @(posedge slow_clk);write_instruction(32'hfc440713); 
    @(posedge slow_clk);write_instruction(32'hfcc40793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'h00c42603); 
    @(posedge slow_clk);write_instruction(32'h01c42583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'ha55ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfc842783); 
    @(posedge slow_clk);write_instruction(32'h02078e63); 
    @(posedge slow_clk);write_instruction(32'h02442703); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f71863); 
    @(posedge slow_clk);write_instruction(32'hfe042703); 
    @(posedge slow_clk);write_instruction(32'h3e700793); 
    @(posedge slow_clk);write_instruction(32'h02e7d263); 
    @(posedge slow_clk);write_instruction(32'hfd840713); 
    @(posedge slow_clk);write_instruction(32'hfc840793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'hfac42603); 
    @(posedge slow_clk);write_instruction(32'h00042583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'ha71ff0ef); 
    @(posedge slow_clk);write_instruction(32'h03c0006f); 
    @(posedge slow_clk);write_instruction(32'hfc842783); 
    @(posedge slow_clk);write_instruction(32'h02078a63); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h02079663); 
    @(posedge slow_clk);write_instruction(32'hfe042703); 
    @(posedge slow_clk);write_instruction(32'h3e700793); 
    @(posedge slow_clk);write_instruction(32'h02e7d063); 
    @(posedge slow_clk);write_instruction(32'hfd840713); 
    @(posedge slow_clk);write_instruction(32'hfc840793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'hfa442603); 
    @(posedge slow_clk);write_instruction(32'h00842583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'ha35ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfc442783); 
    @(posedge slow_clk);write_instruction(32'h02078e63); 
    @(posedge slow_clk);write_instruction(32'h02442703); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'h02f71863); 
    @(posedge slow_clk);write_instruction(32'hfdc42703); 
    @(posedge slow_clk);write_instruction(32'h3e700793); 
    @(posedge slow_clk);write_instruction(32'h02e7d263); 
    @(posedge slow_clk);write_instruction(32'hfd440713); 
    @(posedge slow_clk);write_instruction(32'hfc440793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'hfa842603); 
    @(posedge slow_clk);write_instruction(32'h00442583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'h9f9ff0ef); 
    @(posedge slow_clk);write_instruction(32'h03c0006f); 
    @(posedge slow_clk);write_instruction(32'hfc442783); 
    @(posedge slow_clk);write_instruction(32'h02078a63); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h02079663); 
    @(posedge slow_clk);write_instruction(32'hfdc42703); 
    @(posedge slow_clk);write_instruction(32'h3e700793); 
    @(posedge slow_clk);write_instruction(32'h02e7d063); 
    @(posedge slow_clk);write_instruction(32'hfd440713); 
    @(posedge slow_clk);write_instruction(32'hfc440793); 
    @(posedge slow_clk);write_instruction(32'h00070693); 
    @(posedge slow_clk);write_instruction(32'hfa042603); 
    @(posedge slow_clk);write_instruction(32'h00c42583); 
    @(posedge slow_clk);write_instruction(32'h00078513); 
    @(posedge slow_clk);write_instruction(32'h9bdff0ef); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h02079e63); 
    @(posedge slow_clk);write_instruction(32'hfd442783); 
    @(posedge slow_clk);write_instruction(32'h02078a63); 
    @(posedge slow_clk);write_instruction(32'hfe842783); 
    @(posedge slow_clk);write_instruction(32'h02079663); 
    @(posedge slow_clk);write_instruction(32'hfbc42503); 
    @(posedge slow_clk);write_instruction(32'h909ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00078e63); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hfef42423); 
    @(posedge slow_clk);write_instruction(32'hfac42503); 
    @(posedge slow_clk);write_instruction(32'h8b5ff0ef); 
    @(posedge slow_clk);write_instruction(32'h01042503); 
    @(posedge slow_clk);write_instruction(32'h875ff0ef); 
    @(posedge slow_clk);write_instruction(32'h02442783); 
    @(posedge slow_clk);write_instruction(32'h02079e63); 
    @(posedge slow_clk);write_instruction(32'hfd842783); 
    @(posedge slow_clk);write_instruction(32'h02078a63); 
    @(posedge slow_clk);write_instruction(32'hfe442783); 
    @(posedge slow_clk);write_instruction(32'h02079663); 
    @(posedge slow_clk);write_instruction(32'hfb442503); 
    @(posedge slow_clk);write_instruction(32'h8c9ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00078e63); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hfef42223); 
    @(posedge slow_clk);write_instruction(32'hfa842503); 
    @(posedge slow_clk);write_instruction(32'h875ff0ef); 
    @(posedge slow_clk);write_instruction(32'h01442503); 
    @(posedge slow_clk);write_instruction(32'h835ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00178793); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'hfc842783); 
    @(posedge slow_clk);write_instruction(32'h00078863); 
    @(posedge slow_clk);write_instruction(32'hfe042783); 
    @(posedge slow_clk);write_instruction(32'h00178793); 
    @(posedge slow_clk);write_instruction(32'hfef42023); 
    @(posedge slow_clk);write_instruction(32'hfc442783); 
    @(posedge slow_clk);write_instruction(32'h00078863); 
    @(posedge slow_clk);write_instruction(32'hfdc42783); 
    @(posedge slow_clk);write_instruction(32'h00178793); 
    @(posedge slow_clk);write_instruction(32'hfcf42e23); 
    @(posedge slow_clk);write_instruction(32'hfd842783); 
    @(posedge slow_clk);write_instruction(32'hca0784e3); 
    @(posedge slow_clk);write_instruction(32'hfd442783); 
    @(posedge slow_clk);write_instruction(32'hca0780e3); 
    @(posedge slow_clk);write_instruction(32'h02842783); 
    @(posedge slow_clk);write_instruction(32'hfe842703); 
    @(posedge slow_clk);write_instruction(32'h00e7a023); 
    @(posedge slow_clk);write_instruction(32'h02c42783); 
    @(posedge slow_clk);write_instruction(32'hfe442703); 
    @(posedge slow_clk);write_instruction(32'h00e7a023); 
    @(posedge slow_clk);write_instruction(32'h00000013); 
    @(posedge slow_clk);write_instruction(32'h05c12083); 
    @(posedge slow_clk);write_instruction(32'h05812403); 
    @(posedge slow_clk);write_instruction(32'h06010113); 
    @(posedge slow_clk);write_instruction(32'h00008067); 
    @(posedge slow_clk);write_instruction(32'hf4010113); 
    @(posedge slow_clk);write_instruction(32'h0a112e23); 
    @(posedge slow_clk);write_instruction(32'h0a812c23); 
    @(posedge slow_clk);write_instruction(32'h0a912a23); 
    @(posedge slow_clk);write_instruction(32'h0c010413); 
    @(posedge slow_clk);write_instruction(32'hfe042223); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hfef42023); 
    @(posedge slow_clk);write_instruction(32'h00200793); 
    @(posedge slow_clk);write_instruction(32'hfcf42e23); 
    @(posedge slow_clk);write_instruction(32'h00300793); 
    @(posedge slow_clk);write_instruction(32'hfcf42c23); 
    @(posedge slow_clk);write_instruction(32'h00400793); 
    @(posedge slow_clk);write_instruction(32'hfcf42a23); 
    @(posedge slow_clk);write_instruction(32'h00500793); 
    @(posedge slow_clk);write_instruction(32'hfcf42823); 
    @(posedge slow_clk);write_instruction(32'h00600793); 
    @(posedge slow_clk);write_instruction(32'hfcf42623); 
    @(posedge slow_clk);write_instruction(32'h00700793); 
    @(posedge slow_clk);write_instruction(32'hfcf42423); 
    @(posedge slow_clk);write_instruction(32'h00800793); 
    @(posedge slow_clk);write_instruction(32'hfcf42223); 
    @(posedge slow_clk);write_instruction(32'h00900793); 
    @(posedge slow_clk);write_instruction(32'hfcf42023); 
    @(posedge slow_clk);write_instruction(32'h00a00793); 
    @(posedge slow_clk);write_instruction(32'hfaf42e23); 
    @(posedge slow_clk);write_instruction(32'h00b00793); 
    @(posedge slow_clk);write_instruction(32'hfaf42c23); 
    @(posedge slow_clk);write_instruction(32'h00c00793); 
    @(posedge slow_clk);write_instruction(32'hfaf42a23); 
    @(posedge slow_clk);write_instruction(32'h00d00793); 
    @(posedge slow_clk);write_instruction(32'hfaf42823); 
    @(posedge slow_clk);write_instruction(32'h00e00793); 
    @(posedge slow_clk);write_instruction(32'hfaf42623); 
    @(posedge slow_clk);write_instruction(32'h00f00793); 
    @(posedge slow_clk);write_instruction(32'hfaf42423); 
    @(posedge slow_clk);write_instruction(32'h01000793); 
    @(posedge slow_clk);write_instruction(32'hfaf42223); 
    @(posedge slow_clk);write_instruction(32'h01100793); 
    @(posedge slow_clk);write_instruction(32'hfaf42023); 
    @(posedge slow_clk);write_instruction(32'h01200793); 
    @(posedge slow_clk);write_instruction(32'hf8f42e23); 
    @(posedge slow_clk);write_instruction(32'h01300793); 
    @(posedge slow_clk);write_instruction(32'hf8f42c23); 
    @(posedge slow_clk);write_instruction(32'h01400793); 
    @(posedge slow_clk);write_instruction(32'hf8f42a23); 
    @(posedge slow_clk);write_instruction(32'h01500793); 
    @(posedge slow_clk);write_instruction(32'hf8f42823); 
    @(posedge slow_clk);write_instruction(32'h01600793); 
    @(posedge slow_clk);write_instruction(32'hf8f42623); 
    @(posedge slow_clk);write_instruction(32'h01700793); 
    @(posedge slow_clk);write_instruction(32'hf8f42423); 
    @(posedge slow_clk);write_instruction(32'h01800793); 
    @(posedge slow_clk);write_instruction(32'hf8f42223); 
    @(posedge slow_clk);write_instruction(32'h01900793); 
    @(posedge slow_clk);write_instruction(32'hf8f42023); 
    @(posedge slow_clk);write_instruction(32'h01a00793); 
    @(posedge slow_clk);write_instruction(32'hf6f42e23); 
    @(posedge slow_clk);write_instruction(32'h01b00793); 
    @(posedge slow_clk);write_instruction(32'hf6f42c23); 
    @(posedge slow_clk);write_instruction(32'h01c00793); 
    @(posedge slow_clk);write_instruction(32'hf6f42a23); 
    @(posedge slow_clk);write_instruction(32'h01d00793); 
    @(posedge slow_clk);write_instruction(32'hf6f42823); 
    @(posedge slow_clk);write_instruction(32'h01e00793); 
    @(posedge slow_clk);write_instruction(32'hf6f42623); 
    @(posedge slow_clk);write_instruction(32'h01f00793); 
    @(posedge slow_clk);write_instruction(32'hf6f42423); 
    @(posedge slow_clk);write_instruction(32'hfe042623); 
    @(posedge slow_clk);write_instruction(32'h000f7f13); 
    @(posedge slow_clk);write_instruction(32'hf6042223); 
    @(posedge slow_clk);write_instruction(32'hfc442783); 
    @(posedge slow_clk);write_instruction(32'h00100713); 
    @(posedge slow_clk);write_instruction(32'h00f71733); 
    @(posedge slow_clk);write_instruction(32'hfb442783); 
    @(posedge slow_clk);write_instruction(32'h00100693); 
    @(posedge slow_clk);write_instruction(32'h00f697b3); 
    @(posedge slow_clk);write_instruction(32'h00f76733); 
    @(posedge slow_clk);write_instruction(32'hfc042783); 
    @(posedge slow_clk);write_instruction(32'h00100693); 
    @(posedge slow_clk);write_instruction(32'h00f697b3); 
    @(posedge slow_clk);write_instruction(32'h00f76733); 
    @(posedge slow_clk);write_instruction(32'hfb042783); 
    @(posedge slow_clk);write_instruction(32'h00100693); 
    @(posedge slow_clk);write_instruction(32'h00f697b3); 
    @(posedge slow_clk);write_instruction(32'h00f76733); 
    @(posedge slow_clk);write_instruction(32'hfbc42783); 
    @(posedge slow_clk);write_instruction(32'h00100693); 
    @(posedge slow_clk);write_instruction(32'h00f697b3); 
    @(posedge slow_clk);write_instruction(32'h00f76733); 
    @(posedge slow_clk);write_instruction(32'hfac42783); 
    @(posedge slow_clk);write_instruction(32'h00100693); 
    @(posedge slow_clk);write_instruction(32'h00f697b3); 
    @(posedge slow_clk);write_instruction(32'h00f76733); 
    @(posedge slow_clk);write_instruction(32'hfb842783); 
    @(posedge slow_clk);write_instruction(32'h00100693); 
    @(posedge slow_clk);write_instruction(32'h00f697b3); 
    @(posedge slow_clk);write_instruction(32'h00f76733); 
    @(posedge slow_clk);write_instruction(32'hfa842783); 
    @(posedge slow_clk);write_instruction(32'h00100693); 
    @(posedge slow_clk);write_instruction(32'h00f697b3); 
    @(posedge slow_clk);write_instruction(32'h00f767b3); 
    @(posedge slow_clk);write_instruction(32'hf6442703); 
    @(posedge slow_clk);write_instruction(32'h00f767b3); 
    @(posedge slow_clk);write_instruction(32'hf6f42223); 
    @(posedge slow_clk);write_instruction(32'hf6442783); 
    @(posedge slow_clk);write_instruction(32'h00ff6f33); 
    @(posedge slow_clk);write_instruction(32'hfe042423); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'he80ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050493); 
    @(posedge slow_clk);write_instruction(32'hfe042503); 
    @(posedge slow_clk);write_instruction(32'he74ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00f484b3); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'he64ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00f484b3); 
    @(posedge slow_clk);write_instruction(32'hfd842503); 
    @(posedge slow_clk);write_instruction(32'he54ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00f484b3); 
    @(posedge slow_clk);write_instruction(32'hfd442503); 
    @(posedge slow_clk);write_instruction(32'he44ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00f484b3); 
    @(posedge slow_clk);write_instruction(32'hfd042503); 
    @(posedge slow_clk);write_instruction(32'he34ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00f484b3); 
    @(posedge slow_clk);write_instruction(32'hfcc42503); 
    @(posedge slow_clk);write_instruction(32'he24ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00f484b3); 
    @(posedge slow_clk);write_instruction(32'hfc842503); 
    @(posedge slow_clk);write_instruction(32'he14ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00f487b3); 
    @(posedge slow_clk);write_instruction(32'hf6f42023); 
    @(posedge slow_clk);write_instruction(32'hf6042783); 
    @(posedge slow_clk);write_instruction(32'h54078463); 
    @(posedge slow_clk);write_instruction(32'hfe842783); 
    @(posedge slow_clk);write_instruction(32'h00078c63); 
    @(posedge slow_clk);write_instruction(32'hf8442603); 
    @(posedge slow_clk);write_instruction(32'hfa442583); 
    @(posedge slow_clk);write_instruction(32'hfc442503); 
    @(posedge slow_clk);write_instruction(32'hed4ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfe042423); 
    @(posedge slow_clk);write_instruction(32'hf6042703); 
    @(posedge slow_clk);write_instruction(32'h00400793); 
    @(posedge slow_clk);write_instruction(32'h00f70863); 
    @(posedge slow_clk);write_instruction(32'hf6042703); 
    @(posedge slow_clk);write_instruction(32'h00300793); 
    @(posedge slow_clk);write_instruction(32'h1ef71863); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h06079663); 
    @(posedge slow_clk);write_instruction(32'hf7042783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'hf7442783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'hf8042783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'hf8442783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'hf9042783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'hf9442783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'hfa042783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'hfa442783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfb042883); 
    @(posedge slow_clk);write_instruction(32'hfb442803); 
    @(posedge slow_clk);write_instruction(32'hfc042783); 
    @(posedge slow_clk);write_instruction(32'hfc442703); 
    @(posedge slow_clk);write_instruction(32'hfd042683); 
    @(posedge slow_clk);write_instruction(32'hfe042603); 
    @(posedge slow_clk);write_instruction(32'hfd442583); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'hebcff0ef); 
    @(posedge slow_clk);write_instruction(32'h0680006f); 
    @(posedge slow_clk);write_instruction(32'hf6842783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'hf6c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'hf7842783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'hf7c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'hf8842783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'hf8c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'hf9842783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'hf9c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfa842883); 
    @(posedge slow_clk);write_instruction(32'hfac42803); 
    @(posedge slow_clk);write_instruction(32'hfb842783); 
    @(posedge slow_clk);write_instruction(32'hfbc42703); 
    @(posedge slow_clk);write_instruction(32'hfc842683); 
    @(posedge slow_clk);write_instruction(32'hfd842603); 
    @(posedge slow_clk);write_instruction(32'hfcc42583); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'he54ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00278713); 
    @(posedge slow_clk);write_instruction(32'h41f75793); 
    @(posedge slow_clk);write_instruction(32'h01e7d793); 
    @(posedge slow_clk);write_instruction(32'h00f70733); 
    @(posedge slow_clk);write_instruction(32'h00377713); 
    @(posedge slow_clk);write_instruction(32'h40f707b3); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h06079663); 
    @(posedge slow_clk);write_instruction(32'hf7042783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'hf7442783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'hf8042783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'hf8442783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'hf9042783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'hf9442783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'hfa042783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'hfa442783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfb042883); 
    @(posedge slow_clk);write_instruction(32'hfb442803); 
    @(posedge slow_clk);write_instruction(32'hfc042783); 
    @(posedge slow_clk);write_instruction(32'hfc442703); 
    @(posedge slow_clk);write_instruction(32'hfd042683); 
    @(posedge slow_clk);write_instruction(32'hfe042603); 
    @(posedge slow_clk);write_instruction(32'hfd442583); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'hdc8ff0ef); 
    @(posedge slow_clk);write_instruction(32'h0680006f); 
    @(posedge slow_clk);write_instruction(32'hf6842783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'hf6c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'hf7842783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'hf7c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'hf8842783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'hf8c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'hf9842783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'hf9c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfa842883); 
    @(posedge slow_clk);write_instruction(32'hfac42803); 
    @(posedge slow_clk);write_instruction(32'hfb842783); 
    @(posedge slow_clk);write_instruction(32'hfbc42703); 
    @(posedge slow_clk);write_instruction(32'hfc842683); 
    @(posedge slow_clk);write_instruction(32'hfd842603); 
    @(posedge slow_clk);write_instruction(32'hfcc42583); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'hd60ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00278713); 
    @(posedge slow_clk);write_instruction(32'h41f75793); 
    @(posedge slow_clk);write_instruction(32'h01e7d793); 
    @(posedge slow_clk);write_instruction(32'h00f70733); 
    @(posedge slow_clk);write_instruction(32'h00377713); 
    @(posedge slow_clk);write_instruction(32'h40f707b3); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'h3480006f); 
    @(posedge slow_clk);write_instruction(32'hf6042703); 
    @(posedge slow_clk);write_instruction(32'h00200793); 
    @(posedge slow_clk);write_instruction(32'h00f70863); 
    @(posedge slow_clk);write_instruction(32'hf6042703); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hd4f712e3); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00079a63); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'hbb8ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02079a63); 
    @(posedge slow_clk);write_instruction(32'hfd442503); 
    @(posedge slow_clk);write_instruction(32'hba8ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02079263); 
    @(posedge slow_clk);write_instruction(32'hfe042503); 
    @(posedge slow_clk);write_instruction(32'hb98ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00079a63); 
    @(posedge slow_clk);write_instruction(32'hfd042503); 
    @(posedge slow_clk);write_instruction(32'hb88ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h06078663); 
    @(posedge slow_clk);write_instruction(32'hf7042783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'hf7442783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'hf8042783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'hf8442783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'hf9042783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'hf9442783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'hfa042783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'hfa442783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfb042883); 
    @(posedge slow_clk);write_instruction(32'hfb442803); 
    @(posedge slow_clk);write_instruction(32'hfc042783); 
    @(posedge slow_clk);write_instruction(32'hfc442703); 
    @(posedge slow_clk);write_instruction(32'hfd042683); 
    @(posedge slow_clk);write_instruction(32'hfe042603); 
    @(posedge slow_clk);write_instruction(32'hfd442583); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'hc78ff0ef); 
    @(posedge slow_clk);write_instruction(32'h0a80006f); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'hb10ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02079a63); 
    @(posedge slow_clk);write_instruction(32'hfcc42503); 
    @(posedge slow_clk);write_instruction(32'hb00ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02079263); 
    @(posedge slow_clk);write_instruction(32'hfd842503); 
    @(posedge slow_clk);write_instruction(32'haf0ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00079a63); 
    @(posedge slow_clk);write_instruction(32'hfc842503); 
    @(posedge slow_clk);write_instruction(32'hae0ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h06078463); 
    @(posedge slow_clk);write_instruction(32'hf6842783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'hf6c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'hf7842783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'hf7c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'hf8842783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'hf8c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'hf9842783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'hf9c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfa842883); 
    @(posedge slow_clk);write_instruction(32'hfac42803); 
    @(posedge slow_clk);write_instruction(32'hfb842783); 
    @(posedge slow_clk);write_instruction(32'hfbc42703); 
    @(posedge slow_clk);write_instruction(32'hfc842683); 
    @(posedge slow_clk);write_instruction(32'hfd842603); 
    @(posedge slow_clk);write_instruction(32'hfcc42583); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'hbd0ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00278713); 
    @(posedge slow_clk);write_instruction(32'h41f75793); 
    @(posedge slow_clk);write_instruction(32'h01e7d793); 
    @(posedge slow_clk);write_instruction(32'h00f70733); 
    @(posedge slow_clk);write_instruction(32'h00377713); 
    @(posedge slow_clk);write_instruction(32'h40f707b3); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00079a63); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'ha44ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02079a63); 
    @(posedge slow_clk);write_instruction(32'hfd442503); 
    @(posedge slow_clk);write_instruction(32'ha34ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02079263); 
    @(posedge slow_clk);write_instruction(32'hfe042503); 
    @(posedge slow_clk);write_instruction(32'ha24ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00079a63); 
    @(posedge slow_clk);write_instruction(32'hfd042503); 
    @(posedge slow_clk);write_instruction(32'ha14ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h08078663); 
    @(posedge slow_clk);write_instruction(32'hf7042783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'hf7442783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'hf8042783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'hf8442783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'hf9042783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'hf9442783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'hfa042783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'hfa442783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfb042883); 
    @(posedge slow_clk);write_instruction(32'hfb442803); 
    @(posedge slow_clk);write_instruction(32'hfc042783); 
    @(posedge slow_clk);write_instruction(32'hfc442703); 
    @(posedge slow_clk);write_instruction(32'hfd042683); 
    @(posedge slow_clk);write_instruction(32'hfe042603); 
    @(posedge slow_clk);write_instruction(32'hfd442583); 
    @(posedge slow_clk);write_instruction(32'hfe442503); 
    @(posedge slow_clk);write_instruction(32'hb04ff0ef); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00278713); 
    @(posedge slow_clk);write_instruction(32'h41f75793); 
    @(posedge slow_clk);write_instruction(32'h01e7d793); 
    @(posedge slow_clk);write_instruction(32'h00f70733); 
    @(posedge slow_clk);write_instruction(32'h00377713); 
    @(posedge slow_clk);write_instruction(32'h40f707b3); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'h0ec0006f); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'h97cff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02079a63); 
    @(posedge slow_clk);write_instruction(32'hfcc42503); 
    @(posedge slow_clk);write_instruction(32'h96cff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h02079263); 
    @(posedge slow_clk);write_instruction(32'hfd842503); 
    @(posedge slow_clk);write_instruction(32'h95cff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'h00079a63); 
    @(posedge slow_clk);write_instruction(32'hfc842503); 
    @(posedge slow_clk);write_instruction(32'h94cff0ef); 
    @(posedge slow_clk);write_instruction(32'h00050793); 
    @(posedge slow_clk);write_instruction(32'hac0780e3); 
    @(posedge slow_clk);write_instruction(32'hf6842783); 
    @(posedge slow_clk);write_instruction(32'h00f12e23); 
    @(posedge slow_clk);write_instruction(32'hf6c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12c23); 
    @(posedge slow_clk);write_instruction(32'hf7842783); 
    @(posedge slow_clk);write_instruction(32'h00f12a23); 
    @(posedge slow_clk);write_instruction(32'hf7c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12823); 
    @(posedge slow_clk);write_instruction(32'hf8842783); 
    @(posedge slow_clk);write_instruction(32'h00f12623); 
    @(posedge slow_clk);write_instruction(32'hf8c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12423); 
    @(posedge slow_clk);write_instruction(32'hf9842783); 
    @(posedge slow_clk);write_instruction(32'h00f12223); 
    @(posedge slow_clk);write_instruction(32'hf9c42783); 
    @(posedge slow_clk);write_instruction(32'h00f12023); 
    @(posedge slow_clk);write_instruction(32'hfa842883); 
    @(posedge slow_clk);write_instruction(32'hfac42803); 
    @(posedge slow_clk);write_instruction(32'hfb842783); 
    @(posedge slow_clk);write_instruction(32'hfbc42703); 
    @(posedge slow_clk);write_instruction(32'hfc842683); 
    @(posedge slow_clk);write_instruction(32'hfd842603); 
    @(posedge slow_clk);write_instruction(32'hfcc42583); 
    @(posedge slow_clk);write_instruction(32'hfdc42503); 
    @(posedge slow_clk);write_instruction(32'ha3cff0ef); 
    @(posedge slow_clk);write_instruction(32'hfec42783); 
    @(posedge slow_clk);write_instruction(32'h00278713); 
    @(posedge slow_clk);write_instruction(32'h41f75793); 
    @(posedge slow_clk);write_instruction(32'h01e7d793); 
    @(posedge slow_clk);write_instruction(32'h00f70733); 
    @(posedge slow_clk);write_instruction(32'h00377713); 
    @(posedge slow_clk);write_instruction(32'h40f707b3); 
    @(posedge slow_clk);write_instruction(32'hfef42623); 
    @(posedge slow_clk);write_instruction(32'ha39ff06f); 
    @(posedge slow_clk);write_instruction(32'hfe842783); 
    @(posedge slow_clk);write_instruction(32'ha20798e3); 
    @(posedge slow_clk);write_instruction(32'hfc442503); 
    @(posedge slow_clk);write_instruction(32'h870ff0ef); 
    @(posedge slow_clk);write_instruction(32'hf8442503); 
    @(posedge slow_clk);write_instruction(32'h830ff0ef); 
    @(posedge slow_clk);write_instruction(32'h00100793); 
    @(posedge slow_clk);write_instruction(32'hfef42423); 
    @(posedge slow_clk);write_instruction(32'ha15ff06f); 
    @(posedge slow_clk);write_instruction(32'hffffffff); 
    @(posedge slow_clk);write_instruction(32'hffffffff); 

     $display("Test Results:");
     $display("    PASSES: %d", passes);
     $display("    FAILS : %d", fails);
    #100000
    $display("Finish simulation at time %d", $time);
    $finish;
end

 wrapper dut (
.clk        (clk          ), // Top level system clock input.
.resetn       (resetn       ), // Asynchronous active low reset.
.uart_rxd     (uart_rxd     ), // UART Recieve pin.
.uart_rx_en   (uart_rx_en   ), // Recieve enable
.uart_rx_break(uart_rx_break), // Did we get a BREAK message?
.uart_rx_valid(uart_rx_valid), // Valid data recieved and available.
.uart_rx_data (uart_rx_data ), 
.input_gpio_pins(input_wires), 
.output_gpio_pins(output_wires), 
.write_done(write_done)
); 



endmodule
